-- bring in necessary libraries
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library opcodes;
use opcodes.opcodes.all;

library ALUCommands;
use ALUCommands.ALUCommands.all;

entity AVRControl is
    port (
        );
end AVRControl;

architecture DataFlow of AVRControl is
begin
end DataFlow;



----------------------------------------------------------------------------------
-- Company:         Caltech EE 119B
-- Engineer:        Albert Gural and Bryan He
-- 
-- Design Name:     AVR-Processor
-- Module Name:     Progmem - DataFlow 
-- Project Name:    AVR-Processor
-- Target Devices:  Xilinx Spartan III XC3S1200EFGG3204C
-- Tool versions:   Xilinx ISE 14.7
-- Description:     This component just describes a simple program ROM for the
--                  AVR CPU.
--
-- Revision: 1.0
-- For file history, see https://github.com/agural/AVR-Processor 
--
----------------------------------------------------------------------------------

--
--  PROG_MEMORY
--
--  This is the program memory component.  It is just a fixed ROM with no
--  timing information.  It is meant to be connected to the AVR CPU. The ROM
--  is always enabled and may be changed when Reset it active.
--
--  Inputs:
--    ProgAB - address bus (16 bits)
--    Reset  - system reset (active low)
--
--  Outputs:
--    ProgDB - program memory data bus (16 bits)
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;


entity ProgMemory is
    port (
        ProgAB  :  in   std_logic_vector(15 downto 0);  -- program address bus
        Reset   :  in   std_logic;                      -- system reset
        ProgDB  :  out  std_logic_vector(15 downto 0)   -- program data bus
    );
end ProgMemory;


architecture ROM of ProgMemory is

    -- define the type for the ROM (an array)
    type  ROMtype  is array(0 to 1618) of std_logic_vector(15 downto 0);

    -- define the actual ROM (initialized to a simple program)
    signal  ROMbits  :  ROMtype  :=  (
        X"9488", X"F100", X"94F8", X"F0F7", X"94C8", X"F0E4", X"94B8", X"F0D3", 
        X"9498", X"F0C1", X"94D8", X"F0B5", X"94A8", X"F0A2", X"94E8", X"F096", 
        X"9448", X"F484", X"9418", X"F471", X"9478", X"F467", X"9408", X"F450", 
        X"9428", X"F442", X"9468", X"F436", X"9458", X"F425", X"9438", X"F413", 
        X"940C", X"0025", X"E800", X"940C", X"0651", X"EF0F", X"3F0F", X"F459", 
        X"E000", X"3000", X"F441", X"E505", X"3505", X"F429", X"EA0A", X"3A0A", 
        X"F411", X"940C", X"0036", X"E801", X"940C", X"0651", X"EF0F", X"2E00", 
        X"2E10", X"2E20", X"2E30", X"2E40", X"2E50", X"2E60", X"2E70", X"2E80", 
        X"2E90", X"2EA0", X"2EB0", X"2EC0", X"2ED0", X"2EE0", X"2EF0", X"2F10", 
        X"2F20", X"2F30", X"2F40", X"2F50", X"2F60", X"2F70", X"2F80", X"2F90", 
        X"2FA0", X"2FB0", X"2FC0", X"2FD0", X"2FE0", X"2FF0", X"1500", X"F5F1", 
        X"1501", X"F5E1", X"1502", X"F5D1", X"1503", X"F5C1", X"1504", X"F5B1", 
        X"1505", X"F5A1", X"1506", X"F591", X"1507", X"F581", X"1508", X"F571", 
        X"1509", X"F561", X"150A", X"F551", X"150B", X"F541", X"150C", X"F531", 
        X"150D", X"F521", X"150E", X"F511", X"150F", X"F501", X"1701", X"F4F1", 
        X"1702", X"F4E1", X"1703", X"F4D1", X"1704", X"F4C1", X"1705", X"F4B1", 
        X"1706", X"F4A1", X"1707", X"F491", X"1708", X"F481", X"1709", X"F471", 
        X"170A", X"F461", X"170B", X"F451", X"170C", X"F441", X"170D", X"F431", 
        X"170E", X"F421", X"170F", X"F411", X"940C", X"0099", X"E802", X"940C", 
        X"0651", X"E000", X"2E00", X"2E10", X"2E20", X"2E30", X"2E40", X"2E50", 
        X"2E60", X"2E70", X"2E80", X"2E90", X"2EA0", X"2EB0", X"2EC0", X"2ED0", 
        X"2EE0", X"2EF0", X"2F10", X"2F20", X"2F30", X"2F40", X"2F50", X"2F60", 
        X"2F70", X"2F80", X"2F90", X"2FA0", X"2FB0", X"2FC0", X"2FD0", X"2FE0", 
        X"2FF0", X"1500", X"F5F1", X"1501", X"F5E1", X"1502", X"F5D1", X"1503", 
        X"F5C1", X"1504", X"F5B1", X"1505", X"F5A1", X"1506", X"F591", X"1507", 
        X"F581", X"1508", X"F571", X"1509", X"F561", X"150A", X"F551", X"150B", 
        X"F541", X"150C", X"F531", X"150D", X"F521", X"150E", X"F511", X"150F", 
        X"F501", X"1701", X"F4F1", X"1702", X"F4E1", X"1703", X"F4D1", X"1704", 
        X"F4C1", X"1705", X"F4B1", X"1706", X"F4A1", X"1707", X"F491", X"1708", 
        X"F481", X"1709", X"F471", X"170A", X"F461", X"170B", X"F451", X"170C", 
        X"F441", X"170D", X"F431", X"170E", X"F421", X"170F", X"F411", X"940C", 
        X"00FC", X"E803", X"940C", X"0651", X"9468", X"F947", X"F953", X"F961", 
        X"F976", X"F980", X"F995", X"F9A4", X"F9B2", X"3840", X"F481", X"3058", 
        X"F471", X"3062", X"F461", X"3470", X"F451", X"3081", X"F441", X"3290", 
        X"F431", X"31A0", X"F421", X"30B4", X"F411", X"940C", X"011A", X"E804", 
        X"940C", X"0651", X"ED4F", X"2E84", X"E044", X"2E94", X"E74F", X"2EA4", 
        X"E041", X"2EB4", X"EF4D", X"2EC4", X"E440", X"2ED4", X"EF47", X"2EE4", 
        X"E140", X"2EF4", X"FA85", X"F086", X"FA92", X"F476", X"FAA7", X"F066", 
        X"FAB0", X"F456", X"FAC1", X"F046", X"FAD6", X"F436", X"FAE3", X"F026", 
        X"FAF4", X"F416", X"940C", X"013F", X"E805", X"940C", X"0651", X"EF0F", 
        X"EF1F", X"E020", X"E730", X"E040", X"E75E", X"E76E", X"E870", X"E485", 
        X"E890", X"EFA0", X"EFBF", X"E5C5", X"EADA", X"E7E0", X"E3FF", X"1F01", 
        X"F568", X"F562", X"F55C", X"F555", X"F149", X"F143", X"3F0E", X"F531", 
        X"1F02", X"F522", X"F51C", X"F110", X"F109", X"F103", X"F0FD", X"3F0E", 
        X"F4E9", X"1F21", X"F4DA", X"F4D4", X"F0C8", X"F0C1", X"F0BB", X"F0B5", 
        X"3F2F", X"F4A1", X"1F95", X"F492", X"F48C", X"F080", X"F079", X"F073", 
        X"F06D", X"3F9E", X"F459", X"1D60", X"F048", X"F041", X"F03A", X"F033", 
        X"F02C", X"F025", X"376E", X"F411", X"940C", X"0181", X"E806", X"940C", 
        X"0651", X"0F95", X"F520", X"F119", X"F112", X"F10B", X"F104", X"F4FD", 
        X"379C", X"F4E9", X"0F01", X"F4D8", X"F0D1", X"F4CA", X"F0C3", X"F4BC", 
        X"F4B5", X"3F0D", X"F4A1", X"0F24", X"F090", X"F089", X"F482", X"F07B", 
        X"F474", X"F06D", X"3F2F", X"F459", X"0D70", X"F048", X"F041", X"F43A", 
        X"F033", X"F42C", X"F025", X"3870", X"F411", X"940C", X"01AA", X"E807", 
        X"940C", X"0651", X"9600", X"F0B0", X"F0A9", X"F0A2", X"F09B", X"F094", 
        X"F08D", X"3485", X"F479", X"379C", X"F469", X"9650", X"F458", X"F451", 
        X"F04A", X"F043", X"F03C", X"F035", X"30A0", X"F421", X"30B0", X"F411", 
        X"940C", X"01C5", X"E808", X"940C", X"0651", X"231C", X"F0C8", X"F0C1", 
        X"F0BA", X"F0B3", X"F0AC", X"F0A5", X"3515", X"F491", X"231D", X"F080", 
        X"F479", X"F072", X"F06B", X"F064", X"F05D", X"F451", X"20D0", X"F040", 
        X"F439", X"F032", X"F02B", X"F024", X"F01D", X"F411", X"940C", X"01E3", 
        X"E809", X"940C", X"0651", X"7FCF", X"F1D0", X"F1C9", X"F1C2", X"F1BB", 
        X"F1B4", X"F1AD", X"35C5", X"F599", X"70C0", X"F188", X"F581", X"F17A", 
        X"F173", X"F16C", X"F165", X"30C0", X"F551", X"E5C5", X"EF0F", X"7F0F", 
        X"F130", X"F129", X"F522", X"F11B", X"F514", X"F10D", X"3F0F", X"F4F9", 
        X"7000", X"F0E8", X"F4E1", X"F0DA", X"F0D3", X"F0CC", X"F0C5", X"3000", 
        X"F4B1", X"EF0F", X"7FDF", X"F098", X"F091", X"F48A", X"F083", X"F47C", 
        X"F075", X"3ADA", X"F461", X"70D0", X"F050", X"F449", X"F042", X"F03B", 
        X"F034", X"F02D", X"30D0", X"F419", X"EADA", X"940C", X"0222", X"E80A", 
        X"940C", X"0651", X"9505", X"F4E0", X"F0D9", X"F4D2", X"F0CB", X"F4C4", 
        X"F0BD", X"3F0F", X"F4A9", X"95B5", X"F098", X"F491", X"F08A", X"F083", 
        X"F07C", X"F075", X"30B0", X"F461", X"95E5", X"F050", X"F049", X"F042", 
        X"F03B", X"F034", X"F02D", X"33E8", X"F419", X"9485", X"940C", X"0243", 
        X"E80B", X"940C", X"0651", X"9500", X"F520", X"F519", X"F112", X"F10B", 
        X"F104", X"F0FD", X"3000", X"F4E9", X"9500", X"F4D8", X"F0D1", X"F4CA", 
        X"F0C3", X"F4BC", X"F0B5", X"3F0F", X"F4A1", X"95C0", X"F490", X"F089", 
        X"F482", X"F07B", X"F474", X"F06D", X"3ACA", X"F459", X"95C0", X"F448", 
        X"F041", X"F03A", X"F033", X"F02C", X"F025", X"35C5", X"F411", X"940C", 
        X"026C", X"E80C", X"940C", X"0651", X"1710", X"F4C0", X"F0B9", X"F0B2", 
        X"F0AB", X"F0A4", X"F49D", X"175A", X"F088", X"F081", X"F07A", X"F073", 
        X"F06C", X"F065", X"E400", X"2E30", X"EF0F", X"15F3", X"F438", X"F031", 
        X"F42A", X"F023", X"F41C", X"F015", X"940C", X"0289", X"E80D", X"940C", 
        X"0651", X"0710", X"F4E0", X"F0D9", X"F0D2", X"F0CB", X"F0C4", X"F4BD", 
        X"0751", X"F0A8", X"F0A1", X"F09A", X"F093", X"F08C", X"F085", X"0715", 
        X"F470", X"F069", X"F462", X"F05B", X"F454", X"F44D", X"0750", X"F438", 
        X"F031", X"F02A", X"F023", X"F01C", X"F415", X"940C", X"02AA", X"E80E", 
        X"940C", X"0651", X"E4E0", X"E7FF", X"371F", X"F4A8", X"F0A1", X"F49A", 
        X"F093", X"F48C", X"F485", X"37E0", X"F470", X"F069", X"F462", X"F05B", 
        X"F454", X"F04D", X"3AF0", X"F438", X"F031", X"F42A", X"F423", X"F01C", 
        X"F015", X"940C", X"02C6", X"E80F", X"940C", X"0651", X"2FE3", X"951A", 
        X"F540", X"F139", X"F532", X"F12B", X"F524", X"F11D", X"3F1F", X"F509", 
        X"E800", X"2E00", X"940A", X"F0E8", X"F0E1", X"F0DA", X"F4D3", X"F4CC", 
        X"F0C5", X"2D00", X"370F", X"F4A9", X"EF0F", X"95EA", X"F090", X"F089", 
        X"F082", X"F07B", X"F074", X"F06D", X"36EF", X"F459", X"951A", X"F048", 
        X"F041", X"F43A", X"F033", X"F42C", X"F025", X"3F1E", X"F411", X"940C", 
        X"02F4", X"E900", X"940C", X"0651", X"2F1C", X"271D", X"F170", X"F169", 
        X"F562", X"F15B", X"F554", X"F14D", X"3F1F", X"F539", X"271C", X"F128", 
        X"F121", X"F51A", X"F113", X"F50C", X"F105", X"3A1A", X"F4F1", X"E020", 
        X"2721", X"F0D8", X"F0D1", X"F4CA", X"F0C3", X"F4BC", X"F0B5", X"3A2A", 
        X"F4A1", X"2720", X"F090", X"F089", X"F082", X"F07B", X"F074", X"F06D", 
        X"3525", X"F459", X"2788", X"F048", X"F441", X"F03A", X"F033", X"F02C", 
        X"F025", X"3080", X"F411", X"940C", X"0328", X"E901", X"940C", X"0651", 
        X"9583", X"F138", X"F131", X"F12A", X"F123", X"F11C", X"F115", X"3081", 
        X"F501", X"EF6E", X"9563", X"F0E8", X"F0E1", X"F4DA", X"F0D3", X"F4CC", 
        X"F0C5", X"3F6F", X"F4B1", X"9563", X"F0A0", X"F499", X"F092", X"F08B", 
        X"F084", X"F07D", X"3060", X"F469", X"9403", X"F058", X"F051", X"F44A", 
        X"F443", X"F03C", X"F035", X"2D00", X"3800", X"EF0F", X"F411", X"940C", 
        X"0354", X"E902", X"940C", X"0651", X"95AA", X"E8F0", X"95A6", X"F520", 
        X"F119", X"F112", X"F50B", X"F504", X"F0FD", X"37AF", X"F4E9", X"95E6", 
        X"F4D8", X"F0D1", X"F0CA", X"F4C3", X"F4BC", X"F0B5", X"33E7", X"F4A1", 
        X"9546", X"F090", X"F489", X"F082", X"F07B", X"F074", X"F06D", X"3040", 
        X"F459", X"95F6", X"F048", X"F041", X"F03A", X"F033", X"F02C", X"F025", 
        X"34F0", X"F411", X"940C", X"037F", X"E903", X"940C", X"0651", X"9501", 
        X"F530", X"F129", X"F122", X"F11B", X"F114", X"F50D", X"3001", X"F4F9", 
        X"9561", X"F0E8", X"F4E1", X"F0DA", X"F0D3", X"F0CC", X"F0C5", X"3060", 
        X"F4B1", X"9401", X"F4A0", X"F099", X"F492", X"F48B", X"F084", X"F07D", 
        X"2D00", X"3800", X"EF0F", X"F459", X"9551", X"F448", X"F041", X"F43A", 
        X"F033", X"F42C", X"F425", X"3852", X"F411", X"940C", X"03AA", X"E904", 
        X"940C", X"0651", X"2B21", X"F0D8", X"F0D1", X"F4CA", X"F0C3", X"F4BC", 
        X"F0B5", X"3F2F", X"F4A1", X"2B2C", X"F090", X"F089", X"F482", X"F07B", 
        X"F474", X"F06D", X"3F2F", X"F459", X"2B61", X"F048", X"F041", X"F43A", 
        X"F033", X"F42C", X"F025", X"3A6A", X"F411", X"940C", X"03CA", X"E905", 
        X"940C", X"0651", X"6F1F", X"F090", X"F089", X"F482", X"F07B", X"F474", 
        X"F06D", X"3F1F", X"F459", X"679D", X"F048", X"F041", X"F03A", X"F033", 
        X"F02C", X"F025", X"379D", X"F411", X"940C", X"03E1", X"E906", X"940C", 
        X"0651", X"9408", X"9517", X"F590", X"F189", X"F582", X"F17B", X"F574", 
        X"F16D", X"3F1F", X"F559", X"9408", X"9537", X"F140", X"F139", X"F532", 
        X"F52B", X"F124", X"F11D", X"3B38", X"F509", X"E001", X"9507", X"F4F0", 
        X"F4E9", X"F0E2", X"F4DB", X"F4D4", X"F0CD", X"3000", X"F4B9", X"9408", 
        X"9407", X"F0A0", X"F099", X"F492", X"F48B", X"F084", X"F07D", X"2D00", 
        X"3C00", X"E000", X"F459", X"9507", X"F048", X"F441", X"F03A", X"F033", 
        X"F02C", X"F025", X"3000", X"F411", X"940C", X"0419", X"E907", X"940C", 
        X"0651", X"E5F0", X"0B01", X"F4F8", X"F0F1", X"F0EA", X"F0E3", X"F0DC", 
        X"F4D5", X"3001", X"F4C1", X"9408", X"47F0", X"F4A8", X"F0A1", X"F49A", 
        X"F093", X"F48C", X"F485", X"3DFF", X"F471", X"9408", X"0AA4", X"F058", 
        X"F051", X"F04A", X"F043", X"F03C", X"F035", X"2D0A", X"370E", X"E001", 
        X"F411", X"940C", X"043E", X"E908", X"940C", X"0651", X"E79F", X"E781", 
        X"47AF", X"F0E0", X"F4D9", X"F0D2", X"F0CB", X"F0C4", X"F0BD", X"30A0", 
        X"F4A9", X"0B91", X"F498", X"F091", X"F48A", X"F483", X"F07C", X"F075", 
        X"3890", X"F461", X"9408", X"4A80", X"F448", X"F041", X"F43A", X"F433", 
        X"F02C", X"F025", X"3D80", X"F411", X"940C", X"0461", X"E909", X"940C", 
        X"0651", X"E08D", X"E090", X"9740", X"F4B0", X"F0A9", X"F4A2", X"F09B", 
        X"F494", X"F08D", X"3F8D", X"F479", X"3F9F", X"F469", X"9700", X"F058", 
        X"F051", X"F44A", X"F043", X"F43C", X"F035", X"3F8D", X"F421", X"3F9F", 
        X"F411", X"940C", X"047E", X"E90A", X"940C", X"0651", X"E7EF", X"E7FF", 
        X"1B01", X"F4D8", X"F0D1", X"F0CA", X"F0C3", X"F0BC", X"F4B5", X"3002", 
        X"F4A1", X"1BE1", X"F490", X"F089", X"F482", X"F47B", X"F074", X"F06D", 
        X"38E0", X"F459", X"1BF4", X"F048", X"F041", X"F03A", X"F033", X"F02C", 
        X"F025", X"37FF", X"F411", X"940C", X"04A0", X"E90B", X"940C", X"0651", 
        X"E5E0", X"E7F1", X"574F", X"F4D8", X"F0D1", X"F4CA", X"F0C3", X"F4BC", 
        X"F4B5", X"3841", X"F4A1", X"57E0", X"F490", X"F089", X"F482", X"F07B", 
        X"F474", X"F06D", X"3EE0", X"F459", X"5AF0", X"F448", X"F041", X"F43A", 
        X"F433", X"F02C", X"F025", X"3DF1", X"F411", X"940C", X"04C2", X"E90C", 
        X"940C", X"0651", X"9552", X"F0E8", X"F4E1", X"F0DA", X"F0D3", X"F0CC", 
        X"F0C5", X"3258", X"F4B1", X"94A2", X"F0A0", X"F499", X"F092", X"F08B", 
        X"F084", X"F07D", X"2D0A", X"3E07", X"E002", X"F459", X"95B2", X"F048", 
        X"F441", X"F03A", X"F033", X"F02C", X"F025", X"30B0", X"F411", X"940C", 
        X"04E4", X"E90D", X"940C", X"0651", X"93AF", X"93BF", X"93CF", X"93DF", 
        X"93EF", X"93FF", X"91AF", X"91BF", X"91CF", X"91DF", X"91EF", X"91FF", 
        X"3DA1", X"F461", X"3EB0", X"F451", X"3ACA", X"F441", X"35D5", X"F431", 
        X"30E0", X"F421", X"30F0", X"F411", X"940C", X"0501", X"E90E", X"940C", 
        X"0651", X"EFBF", X"EFAF", X"EFDF", X"ECC0", X"E0F0", X"E8E0", X"E505", 
        X"9300", X"5555", X"EA0A", X"9300", X"AAAA", X"E000", X"9300", X"1234", 
        X"EF0F", X"9300", X"4321", X"E60E", X"9300", X"6E6E", X"9100", X"5555", 
        X"3505", X"F491", X"9100", X"AAAA", X"3A0A", X"F471", X"9100", X"1234", 
        X"3000", X"F451", X"9100", X"4321", X"3F0F", X"F431", X"9100", X"6E6E", 
        X"360E", X"F411", X"940C", X"052F", X"EA00", X"940C", X"0651", X"E021", 
        X"E032", X"E044", X"E150", X"E260", X"E470", X"933C", X"910C", X"3002", 
        X"F511", X"937E", X"910C", X"3400", X"F4F1", X"932D", X"910E", X"3001", 
        X"F4D1", X"910D", X"936D", X"910E", X"3200", X"F4A9", X"910D", X"3200", 
        X"F491", X"935C", X"910C", X"3100", X"F471", X"910E", X"3200", X"F459", 
        X"910E", X"3001", X"F441", X"910D", X"3001", X"F429", X"910D", X"3200", 
        X"F411", X"940C", X"055E", X"EA01", X"940C", X"0651", X"9329", X"9339", 
        X"8348", X"935A", X"9361", X"9371", X"8320", X"9332", X"910A", X"3001", 
        X"F4B9", X"9109", X"3001", X"F4A1", X"9109", X"3100", X"F489", X"8108", 
        X"3004", X"F471", X"9102", X"3200", X"F459", X"9101", X"3200", X"F441", 
        X"9101", X"3002", X"F429", X"8100", X"3001", X"F411", X"940C", X"0583", 
        X"EA02", X"940C", X"0651", X"EFDF", X"ECC0", X"E0F0", X"E8E0", X"AF2C", 
        X"833A", X"8B4E", X"8359", X"8F36", X"8341", X"AF67", X"A370", X"E0D0", 
        X"E8C1", X"EFFF", X"ECE0", X"AD04", X"3001", X"F4B9", X"8102", X"3002", 
        X"F4A1", X"8906", X"3004", X"F489", X"8101", X"3100", X"F471", X"8D0D", 
        X"3002", X"F459", X"8108", X"3004", X"F441", X"AD0E", X"3200", X"F429", 
        X"8D0F", X"3400", X"F411", X"940C", X"05B0", X"EA03", X"940C", X"0651", 
        X"940C", X"05BB", X"EA04", X"940C", X"0651", X"E56A", X"E57A", X"C008", 
        X"EA06", X"940C", X"0651", X"EA85", X"CFF8", X"EA05", X"940C", X"0651", 
        X"ECE6", X"E0F5", X"9409", X"EA07", X"940C", X"0651", X"940E", X"05C8", 
        X"940E", X"0646", X"33B1", X"F531", X"34C1", X"F521", X"35D9", X"F511", 
        X"E0B0", X"E0C0", X"E0D0", X"D072", X"33B1", X"F4E1", X"34C1", X"F4D1", 
        X"35D9", X"F4C1", X"E0B0", X"E0C0", X"E0D0", X"E4E6", X"E0F6", X"9509", 
        X"33B1", X"F481", X"34C1", X"F471", X"35D9", X"F461", X"94F8", X"940E", 
        X"064A", X"3F9F", X"F439", X"37AF", X"F429", X"36E6", X"F419", X"F417", 
        X"940C", X"05F5", X"EA08", X"940C", X"0651", X"E7CF", X"EFBF", X"17CB", 
        X"F018", X"EB00", X"940C", X"0651", X"EB01", X"F084", X"F079", X"F411", 
        X"940C", X"0651", X"EB02", X"E659", X"0F55", X"F445", X"2BBB", X"F012", 
        X"940C", X"0651", X"EB03", X"2BCC", X"F00A", X"F412", X"940C", X"0651", 
        X"EB04", X"2BBB", X"F5F2", X"1BCB", X"F013", X"940C", X"0651", X"EB05", 
        X"95CA", X"F5BB", X"30B1", X"F5AC", X"94F8", X"F19F", X"940E", X"064A", 
        X"F587", X"FBE1", X"F576", X"FBE3", X"F166", X"0FEE", X"F410", X"940C", 
        X"0651", X"EB06", X"0FEE", X"F528", X"F015", X"940C", X"0651", X"EB07", 
        X"1367", X"C01F", X"1367", X"940C", X"0651", X"1368", X"E860", X"FD66", 
        X"EF6F", X"FD63", X"940C", X"0651", X"FD67", X"EA65", X"FF60", X"E060", 
        X"FF65", X"940C", X"0651", X"FF61", X"940C", X"064E", X"E3B1", X"E4C1", 
        X"E5D9", X"9508", X"EF9F", X"E7AF", X"E6E6", X"9518", X"E000", X"940C", 
        X"064E", X"940C", X"0651"
    );



begin
    -- the address has changed - read the new value
    ProgDB <= ROMbits(CONV_INTEGER(ProgAB)) when (CONV_INTEGER(ProgAB) <= ROMbits'high)  else
              X"E0C0";

    -- process to handle Reset
    process(Reset)
    begin
        -- check if Reset is low now
        if  (Reset = '0')  then
            -- reset is active - initialize the ROM (nothing for now)
        end if;
    end process;
end ROM;

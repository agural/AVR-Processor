-- bring in necessary libraries
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library opcodes;
use opcodes.opcodes.all;

library ALUCommands;
use ALUCommands.ALUCommands.all;

entity AVRRegisters is
    port (
        );
end AVRRegisters;

architecture DataFlow of AVRRegisters is
begin
end DataFlow;


